//
module program (
input  [11:0] address,
output [17:0] instruction,
input         enable,
input         clk);
//
//
wire [13:0] address_a;
wire        pipe_a11;
wire [35:0] data_in_a;
wire [35:0] data_out_a_ll;
wire [35:0] data_out_a_lh;
wire [35:0] data_out_a_hl;
wire [35:0] data_out_a_hh;
wire [13:0] address_b;
wire [35:0] data_in_b_ll;
wire [35:0] data_out_b_ll;
wire [35:0] data_in_b_lh;
wire [35:0] data_out_b_lh;
wire [35:0] data_in_b_hl;
wire [35:0] data_out_b_hl;
wire [35:0] data_in_b_hh;
wire [35:0] data_out_b_hh;
wire        enable_b;
wire        clk_b;
wire  [3:0] we_b;
//
//
assign address_a = {address[10:0], 3'b000};
assign data_in_a = 36'b000000000000000000000000000000000000;
//
FD s6_a11_flop ( .D      (address[11]),
                 .Q      (pipe_a11),
                 .C      (clk));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
 s6_4k_mux0_lut( .I0     (data_out_a_ll[0]),
                 .I1     (data_out_a_hl[0]),
                 .I2     (data_out_a_ll[1]),
                 .I3     (data_out_a_hl[1]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[0]),
                 .O6     (instruction[1]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
 s6_4k_mux2_lut( .I0     (data_out_a_ll[2]),
                 .I1     (data_out_a_hl[2]),
                 .I2     (data_out_a_ll[3]),
                 .I3     (data_out_a_hl[3]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[2]),
                 .O6     (instruction[3]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
 s6_4k_mux4_lut( .I0     (data_out_a_ll[4]),
                 .I1     (data_out_a_hl[4]),
                 .I2     (data_out_a_ll[5]),
                 .I3     (data_out_a_hl[5]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[4]),
                 .O6     (instruction[5]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
 s6_4k_mux6_lut( .I0     (data_out_a_ll[6]),
                 .I1     (data_out_a_hl[6]),
                 .I2     (data_out_a_ll[7]),
                 .I3     (data_out_a_hl[7]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[6]),
                 .O6     (instruction[7]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
 s6_4k_mux8_lut( .I0     (data_out_a_ll[32]),
                 .I1     (data_out_a_hl[32]),
                 .I2     (data_out_a_lh[0]),
                 .I3     (data_out_a_hh[0]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[8]),
                 .O6     (instruction[9]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
s6_4k_mux10_lut( .I0     (data_out_a_lh[1]),
                 .I1     (data_out_a_hh[1]),
                 .I2     (data_out_a_lh[2]),
                 .I3     (data_out_a_hh[2]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[10]),
                 .O6     (instruction[11]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
s6_4k_mux12_lut( .I0     (data_out_a_lh[3]),
                 .I1     (data_out_a_hh[3]),
                 .I2     (data_out_a_lh[4]),
                 .I3     (data_out_a_hh[4]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[12]),
                 .O6     (instruction[13]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
s6_4k_mux14_lut( .I0     (data_out_a_lh[5]),
                 .I1     (data_out_a_hh[5]),
                 .I2     (data_out_a_lh[6]),
                 .I3     (data_out_a_hh[6]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[14]),
                 .O6     (instruction[15]));
//
LUT6_2 # (       .INIT   (64'hFF00F0F0CCCCAAAA))
s6_4k_mux16_lut( .I0     (data_out_a_lh[7]),
                 .I1     (data_out_a_hh[7]),
                 .I2     (data_out_a_lh[32]),
                 .I3     (data_out_a_hh[32]),
                 .I4     (pipe_a11),
                 .I5     (1'b1),
                 .O5     (instruction[16]),
                 .O6     (instruction[17]));
//
assign address_b = 14'b00000000000000;
assign data_in_b_ll = {3'h0, data_out_b_ll[32], 24'b000000000000000000000000, data_out_b_ll[7:0]};
assign data_in_b_lh = {3'h0, data_out_b_lh[32], 24'b000000000000000000000000, data_out_b_lh[7:0]};
assign data_in_b_hl = {3'h0, data_out_b_hl[32], 24'b000000000000000000000000, data_out_b_hl[7:0]};
assign data_in_b_hh = {3'h0, data_out_b_hh[32], 24'b000000000000000000000000, data_out_b_hh[7:0]};
assign enable_b = 1'b0;
assign we_b = 4'b0000;
assign clk_b = 1'b0;
//
RAMB16BWER # ( .DATA_WIDTH_A        (9),
               .DOA_REG             (0),
               .EN_RSTRAM_A         ("FALSE"),
               .INIT_A              (32'h000000000),
               .RST_PRIORITY_A      ("CE"),
               .SRVAL_A             (32'h000000000),
               .WRITE_MODE_A        ("WRITE_FIRST"),
               .DATA_WIDTH_B        (9),
               .DOB_REG             (0),
               .EN_RSTRAM_B         ("FALSE"),
               .INIT_B              (32'h000000000),
               .RST_PRIORITY_B      ("CE"),
               .SRVAL_B             (32'h000000000),
               .WRITE_MODE_B        ("WRITE_FIRST"),
               .RSTTYPE             ("SYNC"),
               .INIT_FILE           ("NONE"),
               .SIM_COLLISION_CHECK ("ALL"),
               .SIM_DEVICE          ("SPARTAN6"),
               .INIT_00             (256'h6B656B036B6D6B036B6F6B036B636B036B6C6B036B656B036B776B036B026B00),
               .INIT_01             (256'h6B706B036B6F6B036B6F6B036B4C6B036B206B036B6F6B036B746B036B206B03),
               .INIT_02             (256'h00005E036B036B036B216B036B6B6B036B636B036B616B036B626B036B2D6B03),
               .INIT_03             (256'h0000000000000000000000000000000000006B0E055E036B025E0E04006301FF),
               .INIT_04             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_05             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_06             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_07             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_08             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_09             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_10             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_11             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_12             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_13             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_14             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_15             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_16             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_17             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_18             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_19             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_20             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_21             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_22             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_23             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_24             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_25             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_26             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_27             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_28             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_29             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_30             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_31             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_32             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_33             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_34             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_35             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_36             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_37             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_38             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_39             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_00            (256'h0000000000000000000000000000000000001833955555555555555555555554),
               .INITP_01            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_02            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_03            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_04            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_05            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_06            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_07            (256'h0000000000000000000000000000000000000000000000000000000000000000))
kcpsm6_rom_ll( .ADDRA               (address_a),
               .ENA                 (enable),
               .CLKA                (clk),
               .DOA                 (data_out_a_ll[31:0]),
               .DOPA                (data_out_a_ll[35:32]), 
               .DIA                 (data_in_a[31:0]),
               .DIPA                (data_in_a[35:32]), 
               .WEA                 (4'h0),
               .REGCEA              (1'b0),
               .RSTA                (1'b0),
               .ADDRB               (address_b),
               .ENB                 (enable_b),
               .CLKB                (clk_b),
               .DOB                 (data_out_b_ll[31:0]),
               .DOPB                (data_out_b_ll[35:32]), 
               .DIB                 (data_in_b_ll[31:0]),
               .DIPB                (data_in_b_ll[35:32]), 
               .WEB                 (we_b),
               .REGCEB              (1'b0),
               .RSTB                (1'b0));
//
RAMB16BWER # ( .DATA_WIDTH_A        (9),
               .DOA_REG             (0),
               .EN_RSTRAM_A         ("FALSE"),
               .INIT_A              (32'h000000000),
               .RST_PRIORITY_A      ("CE"),
               .SRVAL_A             (32'h000000000),
               .WRITE_MODE_A        ("WRITE_FIRST"),
               .DATA_WIDTH_B        (9),
               .DOB_REG             (0),
               .EN_RSTRAM_B         ("FALSE"),
               .INIT_B              (32'h000000000),
               .RST_PRIORITY_B      ("CE"),
               .SRVAL_B             (32'h000000000),
               .WRITE_MODE_B        ("WRITE_FIRST"),
               .RSTTYPE             ("SYNC"),
               .INIT_FILE           ("NONE"),
               .SIM_COLLISION_CHECK ("ALL"),
               .SIM_DEVICE          ("SPARTAN6"),
               .INIT_00             (256'h0008006800080068000800680008006800080068000800680008006800080000),
               .INIT_01             (256'h0008006800080068000800680008006800080068000800680008006800080068),
               .INIT_02             (256'h4800106800080068000800680008006800080068000800680008006800080068),
               .INIT_03             (256'h000000000000000000000000000000000028D0A74F10690049F0A04800106838),
               .INIT_04             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_05             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_06             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_07             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_08             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_09             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_10             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_11             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_12             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_13             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_14             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_15             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_16             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_17             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_18             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_19             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_20             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_21             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_22             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_23             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_24             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_25             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_26             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_27             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_28             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_29             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_30             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_31             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_32             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_33             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_34             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_35             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_36             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_37             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_38             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_39             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_00            (256'h00000000000000000000000000000000000067463BBBBBBBBBBBBBBBBBBBBBBA),
               .INITP_01            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_02            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_03            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_04            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_05            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_06            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_07            (256'h0000000000000000000000000000000000000000000000000000000000000000))
kcpsm6_rom_lh( .ADDRA               (address_a),
               .ENA                 (enable),
               .CLKA                (clk),
               .DOA                 (data_out_a_lh[31:0]),
               .DOPA                (data_out_a_lh[35:32]), 
               .DIA                 (data_in_a[31:0]),
               .DIPA                (data_in_a[35:32]), 
               .WEA                 (4'h0),
               .REGCEA              (1'b0),
               .RSTA                (1'b0),
               .ADDRB               (address_b),
               .ENB                 (enable_b),
               .CLKB                (clk_b),
               .DOB                 (data_out_b_lh[31:0]),
               .DOPB                (data_out_b_lh[35:32]), 
               .DIB                 (data_in_b_lh[31:0]),
               .DIPB                (data_in_b_lh[35:32]), 
               .WEB                 (we_b),
               .REGCEB              (1'b0),
               .RSTB                (1'b0));
//
RAMB16BWER # ( .DATA_WIDTH_A        (9),
               .DOA_REG             (0),
               .EN_RSTRAM_A         ("FALSE"),
               .INIT_A              (32'h000000000),
               .RST_PRIORITY_A      ("CE"),
               .SRVAL_A             (32'h000000000),
               .WRITE_MODE_A        ("WRITE_FIRST"),
               .DATA_WIDTH_B        (9),
               .DOB_REG             (0),
               .EN_RSTRAM_B         ("FALSE"),
               .INIT_B              (32'h000000000),
               .RST_PRIORITY_B      ("CE"),
               .SRVAL_B             (32'h000000000),
               .WRITE_MODE_B        ("WRITE_FIRST"),
               .RSTTYPE             ("SYNC"),
               .INIT_FILE           ("NONE"),
               .SIM_COLLISION_CHECK ("ALL"),
               .SIM_DEVICE          ("SPARTAN6"),
               .INIT_00             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_01             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_02             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_03             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_04             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_05             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_06             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_07             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_08             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_09             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_10             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_11             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_12             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_13             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_14             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_15             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_16             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_17             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_18             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_19             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_20             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_21             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_22             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_23             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_24             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_25             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_26             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_27             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_28             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_29             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_30             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_31             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_32             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_33             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_34             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_35             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_36             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_37             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_38             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_39             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_00            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_01            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_02            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_03            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_04            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_05            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_06            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_07            (256'h0000000000000000000000000000000000000000000000000000000000000000))
kcpsm6_rom_hl( .ADDRA               (address_a),
               .ENA                 (enable),
               .CLKA                (clk),
               .DOA                 (data_out_a_hl[31:0]),
               .DOPA                (data_out_a_hl[35:32]), 
               .DIA                 (data_in_a[31:0]),
               .DIPA                (data_in_a[35:32]), 
               .WEA                 (4'h0),
               .REGCEA              (1'b0),
               .RSTA                (1'b0),
               .ADDRB               (address_b),
               .ENB                 (enable_b),
               .CLKB                (clk_b),
               .DOB                 (data_out_b_hl[31:0]),
               .DOPB                (data_out_b_hl[35:32]), 
               .DIB                 (data_in_b_hl[31:0]),
               .DIPB                (data_in_b_hl[35:32]), 
               .WEB                 (we_b),
               .REGCEB              (1'b0),
               .RSTB                (1'b0));
//
RAMB16BWER # ( .DATA_WIDTH_A        (9),
               .DOA_REG             (0),
               .EN_RSTRAM_A         ("FALSE"),
               .INIT_A              (32'h000000000),
               .RST_PRIORITY_A      ("CE"),
               .SRVAL_A             (32'h000000000),
               .WRITE_MODE_A        ("WRITE_FIRST"),
               .DATA_WIDTH_B        (9),
               .DOB_REG             (0),
               .EN_RSTRAM_B         ("FALSE"),
               .INIT_B              (32'h000000000),
               .RST_PRIORITY_B      ("CE"),
               .SRVAL_B             (32'h000000000),
               .WRITE_MODE_B        ("WRITE_FIRST"),
               .RSTTYPE             ("SYNC"),
               .INIT_FILE           ("NONE"),
               .SIM_COLLISION_CHECK ("ALL"),
               .SIM_DEVICE          ("SPARTAN6"),
               .INIT_00             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_01             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_02             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_03             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_04             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_05             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_06             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_07             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_08             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_09             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_0F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_10             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_11             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_12             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_13             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_14             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_15             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_16             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_17             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_18             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_19             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_1F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_20             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_21             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_22             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_23             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_24             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_25             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_26             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_27             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_28             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_29             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_2F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_30             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_31             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_32             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_33             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_34             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_35             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_36             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_37             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_38             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_39             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3A             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3B             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3C             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3D             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3E             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INIT_3F             (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_00            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_01            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_02            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_03            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_04            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_05            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_06            (256'h0000000000000000000000000000000000000000000000000000000000000000),
               .INITP_07            (256'h0000000000000000000000000000000000000000000000000000000000000000))
kcpsm6_rom_hh( .ADDRA               (address_a),
               .ENA                 (enable),
               .CLKA                (clk),
               .DOA                 (data_out_a_hh[31:0]),
               .DOPA                (data_out_a_hh[35:32]), 
               .DIA                 (data_in_a[31:0]),
               .DIPA                (data_in_a[35:32]), 
               .WEA                 (4'h0),
               .REGCEA              (1'b0),
               .RSTA                (1'b0),
               .ADDRB               (address_b),
               .ENB                 (enable_b),
               .CLKB                (clk_b),
               .DOB                 (data_out_b_hh[31:0]),
               .DOPB                (data_out_b_hh[35:32]), 
               .DIB                 (data_in_b_hh[31:0]),
               .DIPB                (data_in_b_hh[35:32]), 
               .WEB                 (we_b),
               .REGCEB              (1'b0),
               .RSTB                (1'b0));
//
endmodule
